----------------------------------------------------------------------------------
-- Company: FER
-- Engineer: Mrkovic, Ramljak
-- 
-- Create Date: 05/10/2021 04:25:36 PM
-- Design Name: AXI_Network_Adapter
-- Module Name: SNA_resp_buffer_controller - Behavioral
-- Project Name: NoC_Router
-- Target Devices: zc706
-- Tool Versions: 2020.2
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- Revision 0.1 - 2021-05-10 - Ramljak
-- Additional Comments: Prva verzija SNA_resp_buffer_controllera
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

library noc_lib;
use noc_lib.router_config.ALL;
use noc_lib.AXI_network_adapter_config.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
-- use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
-- library UNISIM;
-- use UNISIM.VComponents.all;

entity SNA_resp_buffer_controller is

    Generic (
        flit_size : integer := const_flit_size;
        vc_num : integer := const_vc_num;
        mesh_size_x : integer := const_mesh_size_x;
        mesh_size_y : integer := const_mesh_size_y;
        address_size : integer := const_address_size;
        injection_vc : integer := const_default_injection_vc
    );
                  
    Port (
        clk : in std_logic;
        rst : in std_logic; 
                   
        flit_in : out std_logic_vector(flit_size - 1 downto 0);
        flit_in_valid : out std_logic;
        
        op_write : in std_logic;
        op_read : in std_logic;
        
        data : in std_logic_vector(31 downto 0);
        resp : in std_logic_vector(1 downto 0);
        
        r_addr : in std_logic_vector(address_size - 1 downto 0);
        t_end : out std_logic
    );

end SNA_resp_buffer_controller;

architecture Behavioral of SNA_resp_buffer_controller is

    -- ENUMERACIJA STANJA fsm-a
    type state_type is (IDLE, W_FLIT_1, R_FLIT_1, R_FLIT_2);
    -- TRENUTNO STANJE
    signal current_state : state_type;
    -- SLJEDECE STANJE
    signal next_state : state_type;
    -- POCETNO STANJE
    constant initial_state : state_type := IDLE;

    -- enable SIGNALI PROCESA INDIVIDUALNIH STANJA
    signal W_FLIT_1_enable : std_logic;
    signal R_FLIT_1_enable : std_logic;
    signal R_FLIT_2_enable : std_logic;
begin

    -- PROCES KOJI KOORDINIRA PROCESE POJEDINIH STANJA
    combinatorial_process : process (current_state, op_write, op_read) is
    
    begin
    
        W_FLIT_1_enable <= '0';
        R_FLIT_1_enable <= '0';
        R_FLIT_2_enable <= '0';
        
        t_end <= '0';
    
        case current_state is
        
            when IDLE =>
            
                if op_write = '1' then
                    
                    next_state <= W_FLIT_1;
                    W_FLIT_1_enable <= '1';
                
                elsif op_read = '1' then
                    
                    next_state <= R_FLIT_1;
                    R_FLIT_1_enable <= '1';
                    
                else
                
                    next_state <= IDLE;
                
                end if;   
            
            when W_FLIT_1 =>
            
                next_state <= IDLE;
                
                t_end <= '1';
                
            when R_FLIT_1 =>
            
                next_state <= R_FLIT_2;
                R_FLIT_2_enable <= '1';
                
            when R_FLIT_2 =>
            
                next_state <= IDLE;
                
                t_end <= '1';
            
        end case;
    
    end process;
    
    -- PROCES KOJI GRADI I ODASILJE FLITOVE
    builder_process : process (clk) is
    
        variable flit_var : std_logic_vector(flit_size - 1 downto 0);
        variable flit_valid_var : std_logic;
        variable vc_var : std_logic_vector(vc_num - 1 downto 0);
    
    begin
    
        if rising_edge(clk) then
            if rst = '0' then
                
                -- Varijable
                flit_var := (others => '0');
                flit_valid_var := '0';
                vc_var := (others => '0');
                
                -- Izlazni signali
                flit_in <= (others => '0');
                flit_in_valid <= '0';
                
            else
            
                flit_var := (others => '0');
                flit_valid_var := '0';
                vc_var := (injection_vc => '1', others => '0');
                
                if W_FLIT_1_enable = '1' then
                
                    -- FLIT LABELA
                    flit_var(flit_size - 1 downto flit_size - 2) := "11";
                    -- VIRTUALNI KANAL
                    flit_var(flit_size - 2 - 1 downto flit_size - 2 - vc_num) := vc_var;
                    -- X KOORDNIATA DESTINACIJE
                    flit_var(flit_size - 2 - vc_num - 1 downto
                             flit_size - 2 - vc_num - mesh_size_x) := r_addr(address_size - 1 downto address_size - mesh_size_x); 
                    -- Y KOORDINATA DESTINACIJE
                    flit_var(flit_size - 2 - vc_num - mesh_size_x - 1 downto
                             flit_size - 2 - vc_num - mesh_size_x - mesh_size_y) := r_addr(address_size - mesh_size_x - 1 downto 0);
                    -- WRITE RESPONSE
                    flit_var(2 downto 1) := resp;
                    -- R/W
                    flit_var(0) := '0';
                    
                    flit_valid_var := '1';
                
                elsif R_FLIT_1_enable = '1' then
                
                    -- FLIT LABELA
                    flit_var(flit_size - 1 downto
                             flit_size - 2) := "10";
                    -- VIRTUALNI KANAL
                    flit_var(flit_size - 2 - 1 downto
                             flit_size - 2 - vc_num) := vc_var;
                    -- X KOORDNIATA DESTINACIJE
                    flit_var(flit_size - 2 - vc_num - 1 downto
                             flit_size - 2 - vc_num - mesh_size_x) := r_addr(address_size - 1 downto address_size - mesh_size_x); 
                    -- Y KOORDINATA DESTINACIJE
                    flit_var(flit_size - 2 - vc_num - mesh_size_x - 1 downto
                             flit_size - 2 - vc_num - mesh_size_x - mesh_size_y) := r_addr(address_size - mesh_size_x - 1 downto 0);
                    -- READ RESPONSE
                    flit_var(2 downto 1) := resp;
                    -- R/W
                    flit_var(0) := '1';
                    
                    flit_valid_var := '1';
                
                elsif R_FLIT_2_enable = '1' then
                
                    -- FLIT LABELA
                    flit_var(flit_size - 1 downto
                             flit_size - 2) := "01";
                    -- VIRTUALNI KANAL
                    flit_var(flit_size - 2 - 1 downto
                             flit_size - 2 - vc_num) := vc_var;
                    -- X KOORDNIATA DESTINACIJE
                    flit_var(flit_size - 2 - vc_num - 1 downto
                             flit_size - 2 - vc_num - mesh_size_x) := r_addr(address_size - 1 downto address_size - mesh_size_x); 
                    -- Y KOORDINATA DESTINACIJE
                    flit_var(flit_size - 2 - vc_num - mesh_size_x - 1 downto
                             flit_size - 2 - vc_num - mesh_size_x - mesh_size_y) := r_addr(address_size - mesh_size_x - 1 downto 0);
                    -- READ ADDRESS
                    flit_var(31 downto 0) := data;
                    
                    flit_valid_var := '1';
                
                end if;
                
                flit_in <= flit_var;
                flit_in_valid <= flit_valid_var;
                
            end if;
        end if;
    
    end process;
    
    -- PROCES KOJI IZRACUNAVA TRENUTNO STANJE
    synchronous_process : process (clk) is
    
    begin
        
        if rising_edge(clk) then
            if rst = '0' then
                current_state <= initial_state;
            else
                current_state <= next_state;
            end if;
        end if;    
        
    end process;

end Behavioral;
